//Jack Gentsch, Jacky Wang, Chinh Bui
//Lab 5: Instruction memory module for the cpu
//EE 469 with James Peckol 5/25/16
//A 32 bit wide, 128 words long instruction memory for the cpu
module imem (dataOut, adrx, clk, reset, altProgram);
	output [31:0] dataOut;
	input [6:0] adrx;
	input clk, reset, altProgram;
	
	reg [31:0] mem [0:127];
	
	//Initialization of instructions in memory
	always @(posedge clk) begin
		if (reset) begin
			//if (~altProgram) begin
				$readmemb("mips2mach.txt", mem);
				/*
				mem[0] = 100011_00000_01001_0000000000000000;
				mem[1] = 100011_00000_01010_0000000000000001;
				mem[2] = 001000_00000_01011_0000000000000011;
				mem[3] = 000000_01001_01010_01001_00000_100010;
				mem[4] = 000000_01011_01001_01010_00000_101010;
				mem[5] = 000101_01010_00000_0000000001001000;
				mem[6] = 000000_00000_00000_0000000000000000;

				mem[7] = 100011_00000_01001_0000000000000010;
				mem[8] = 000000_00000_01001_01001_00101_000000;
				mem[9] = 101011_00000_01001_0000000000000010;
				mem[10] = 001000_00000_01100_0000000000000111;
				mem[11] = 101011_00000_01100_0000000000000011;
				mem[12] = 100011_00000_01001_0000000000000100;
				mem[13] = 100011_00000_01010_0000000000000101;
				mem[14] = 000000_01001_01010_01011_00000_100100;
				mem[15] = 101011_00000_01011_0000000000000110;
				mem[16] = 000010_00000000000000000001110100;
				mem[17] = 000000_00000_00000_0000000000000000;

				mem[18] = 100011_00000_01001_0000000000000010;
				mem[19] = 001000_00000_01010_0000000000000100;
				mem[20] = 000000_01001_01010_01001_00000_100000;
				mem[21] = 101011_00000_01001_0000000000000010;
				mem[22] = 001000_00000_01010_0000000000000011;
				mem[23] = 000000_01001_01010_01011_00000_100010;
				mem[24] = 101011_00000_01011_0000000000000011;
				mem[25] = 100011_00000_01001_0000000000000100;
				mem[26] = 100011_00000_01010_0000000000000101;
				mem[27] = 000000_01001_01010_01011_00000_100101;
				mem[28] = 101011_00000_01011_0000000000000110;

				mem[29] = 100011_00000_01001_0000000000000000;
				mem[30] = 100011_00000_01010_0000000000000001;
				mem[31] = 000000_01001_01010_01001_00000_100000;
				mem[32] = 101011_00000_01001_0000000000000000;
				mem[33] = 100011_00000_01001_0000000000000100;
				mem[34] = 100011_00000_01010_0000000000000101;
				mem[35] = 100011_00000_01011_0000000000000111;
				mem[36] = 000000_01001_01010_01001_00000_100110;
				mem[37] = 000000_01001_01001_01011_00000_100100;
				mem[38] = 101011_00000_01001_0000000000000110;
				*/

				// instruction from lab 4
				/*mem[0] = 32'b100011_00000_01001_0000000000000000;
				mem[1] = 32'b100011_00000_01010_0000000000000001;
				mem[2] = 32'b000000_01001_01010_01001_00000_100010;
				mem[3] = 32'b001000_00000_01011_0000000000000011;
				mem[4] = 32'b000000_01011_01001_01010_00000_101010;
				mem[5] = 32'b000101_01010_00000_0000000000110000;
				mem[6] = 32'b100011_00000_01001_0000000000000010;
				mem[7] = 32'b000000_00000_01001_01001_00101_000000;
				mem[8] = 32'b101011_00000_01001_0000000000000010;
				mem[9] = 32'b001000_00000_01100_0000000000000111;
				mem[10] = 32'b101011_00000_01100_0000000000000011;
				mem[11] = 32'b000010_00000000000000000001000100;
				mem[12] = 32'b001000_00000_01100_0000000000000110;
				mem[13] = 32'b101011_00000_01100_0000000000000010;
				mem[14] = 32'b100011_00000_01001_0000000000000011;
				mem[15] = 32'b000000_00000_01001_01001_00010_000000;
				mem[16] = 32'b101011_00000_01001_0000000000000011;
				mem[17] = 32'b111111_00000000000000000000000000;
			end else begin
				mem[0] = 32'b100011_00000_01001_0000000000000000;
				mem[1] = 32'b100011_00000_01010_0000000000000001;
				mem[2] = 32'b000000_01001_01010_01011_00000_100100; //AND 7, 5
				mem[3] = 32'b000000_01001_01010_01000_00000_100101; //OR 7, 5
				mem[4] = 32'b000000_01001_01010_01000_00000_100110; //XOR 7, 5
				mem[5] = 32'b000000_01011_00000_00000_00000_001000; //JR [AND RESULT] == 2 (should loop forever)
				mem[6] = 32'b111111_00000000000000000000000000; //HALT*/
			//end
		end
	end

	assign dataOut = mem[adrx];

endmodule
