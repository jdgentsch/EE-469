// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 14.0.0 Build 200 06/17/2014 SJ Web Edition"
// CREATED		"Wed Oct 14 14:20:43 2015"


/*
IMPORTANT NOTE TO THE GRADER:
This file was generated using a schematic level file, "syncSchematic.bsf"
The file should be attached within our submitted zip file.

Note that the output bus, [3:0]q, were manually assigned on line 73. This was code
written by students, not generated by Quartus. This was according to professor
Peckol's recommendation, as other students have found similar bugs with the 
Verilog synthesizer.

Jack Gentsch and Jacky Wang
10/14/2015
*/

module syncSchematic(
	clk,
	reset,
	q
);


input wire	clk;
input wire	reset;
output wire	[3:0] q;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
reg	SYNTHESIZED_WIRE_15;
reg	SYNTHESIZED_WIRE_16;
reg	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
reg	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;

assign	SYNTHESIZED_WIRE_1 = 1;
assign	SYNTHESIZED_WIRE_3 = 1;
assign	SYNTHESIZED_WIRE_12 = 1;
assign	SYNTHESIZED_WIRE_14 = 1;

//Note these four lines were written by the students
//Read foreword for more information
assign q[3] = SYNTHESIZED_WIRE_18;
assign q[2] = SYNTHESIZED_WIRE_17;
assign q[1] = SYNTHESIZED_WIRE_15;
assign q[0] = SYNTHESIZED_WIRE_16;



always@(posedge clk or negedge reset or negedge SYNTHESIZED_WIRE_1)
begin
if (!reset)
	begin
	SYNTHESIZED_WIRE_16 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_1)
	begin
	SYNTHESIZED_WIRE_16 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_0;
	end
end


always@(posedge clk or negedge reset or negedge SYNTHESIZED_WIRE_3)
begin
if (!reset)
	begin
	SYNTHESIZED_WIRE_15 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_3)
	begin
	SYNTHESIZED_WIRE_15 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_2;
	end
end

assign	SYNTHESIZED_WIRE_2 = SYNTHESIZED_WIRE_15 ~^ SYNTHESIZED_WIRE_16;

assign	SYNTHESIZED_WIRE_5 = SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_16;

assign	SYNTHESIZED_WIRE_4 = SYNTHESIZED_WIRE_17 & SYNTHESIZED_WIRE_15;

assign	SYNTHESIZED_WIRE_0 =  ~SYNTHESIZED_WIRE_16;

assign	SYNTHESIZED_WIRE_6 = ~(SYNTHESIZED_WIRE_17 | SYNTHESIZED_WIRE_15 | SYNTHESIZED_WIRE_16);

assign	SYNTHESIZED_WIRE_11 = SYNTHESIZED_WIRE_4 | SYNTHESIZED_WIRE_5 | SYNTHESIZED_WIRE_6;

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_7 | SYNTHESIZED_WIRE_8 | SYNTHESIZED_WIRE_9 | SYNTHESIZED_WIRE_10;

assign	SYNTHESIZED_WIRE_7 = ~(SYNTHESIZED_WIRE_18 | SYNTHESIZED_WIRE_15 | SYNTHESIZED_WIRE_17 | SYNTHESIZED_WIRE_16);

assign	SYNTHESIZED_WIRE_10 = SYNTHESIZED_WIRE_18 & SYNTHESIZED_WIRE_17;

assign	SYNTHESIZED_WIRE_8 = SYNTHESIZED_WIRE_18 & SYNTHESIZED_WIRE_15;


always@(posedge clk or negedge reset or negedge SYNTHESIZED_WIRE_12)
begin
if (!reset)
	begin
	SYNTHESIZED_WIRE_17 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_12)
	begin
	SYNTHESIZED_WIRE_17 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_11;
	end
end

assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_18 & SYNTHESIZED_WIRE_16;


always@(posedge clk or negedge reset or negedge SYNTHESIZED_WIRE_14)
begin
if (!reset)
	begin
	SYNTHESIZED_WIRE_18 <= 0;
	end
else
if (!SYNTHESIZED_WIRE_14)
	begin
	SYNTHESIZED_WIRE_18 <= 1;
	end
else
	begin
	SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_13;
	end
end






endmodule
