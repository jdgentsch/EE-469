module memoryManager ();
	sram mySRAM ();
	registerFile myRegFile ();

endmodule