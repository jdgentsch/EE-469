//Jack Gentsch, Jacky Wang, Chinh Bui
//Lab 3: ALU
//EE 469 with James Peckol 4/22/16

module alu (out, zero, overflow, cout, neg, busA, busB, control);
	output [31:0] out;
	output zero, overflow, cout, neg;
	input [31:0] busA, busB;
	input [2:0] control;

	

endmodule
