module registerFile ();
	



endmodule