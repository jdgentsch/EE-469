//Jack Gentsch, Jacky Wang, Chinh Bui
//EE 469, Dr. Peckol 4/15/16
// 4-bit Carry Look Ahead (cla) Adder

module cla4 (sum, Cout, pOut, gOut, inA, inB, Cin);
	output [3:0] sum;
	output Cout, pOut, gOut; // pOut = propagate, gOut = generate
	input [3:0] inA, inB;
	input Cin;



endmodule
