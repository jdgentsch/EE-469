//Jack Gentsch, Jacky Wang, Chinh Bui
//Lab 3: ALU with dataflow model
//EE 469 with James Peckol 4/22/16

module alu (busOut, zero, overflow, Cout, neg, busA, busB, control);
	output [31:0] busOut;
	output zero, overflow, Cout, neg;
	input [31:0] busA, busB;
	input [2:0] control;



endmodule
